module BranchPredict();

endmodule