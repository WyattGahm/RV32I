module Registers(input wire [4:0] read1, input wire [4:0] read2, input wire [4:0] write, input wire [31:0] write_data, input wire [0:0] RegWrite, output wire [31:0] out1, output wire [31:0] out2);
	reg [31:0] registers [31:0];
	
	assign out1 = (read1 == 5'd0) ? 32'd0 : registers[read1];
	assign out2 = (read2 == 5'd0) ? 32'd0 : registers[read2];
	
	
	always@(*) begin
		if(RegWrite == 1'b1) registers[write] = write_data; 
	end
	
	
	
	initial begin
		registers[0]  = 32'd0;
		registers[1]  = 32'd0;
		registers[2]  = 32'd0;
		registers[3]  = 32'd0;
		registers[4]  = 32'd0;
		registers[5]  = 32'd0;
		registers[6]  = 32'd0;
		registers[7]  = 32'd0;
		registers[8]  = 32'd0;
		registers[9]  = 32'd0;
		registers[10] = 32'd0;
		registers[11] = 32'd0;
		registers[12] = 32'd0;
		registers[13] = 32'd0;
		registers[14] = 32'd0;
		registers[15] = 32'd0;
		registers[16] = 32'd0;
		registers[17] = 32'd0;
		registers[18] = 32'd0;
		registers[19] = 32'd0;
		registers[20] = 32'd0;
		registers[21] = 32'd0;
		registers[22] = 32'd0;
		registers[23] = 32'd0;
		registers[24] = 32'd0;
		registers[25] = 32'd0;
		registers[26] = 32'd0;
		registers[27] = 32'd0;
		registers[28] = 32'd0;
		registers[29] = 32'd0;
		registers[30] = 32'd0;
		registers[31] = 32'd0;
	end
endmodule